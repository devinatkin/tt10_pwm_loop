/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

`timescale 1ns/1ps

module tt_um_devinatkin_pwm (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output reg  [7:0] uo_out,   // Dedicated outputs
    input  wire       clk,      // Clock
    input  wire       rst_n     // Active-low reset
);

    parameter WIDTH = 8;        // Width of each register
    parameter SIZE = 8;         // Number of registers

    wire slow_clk;  // Slow clock generated by PWM
    reg gated_slow_clk; // Gated slow clock

    wire [WIDTH-1:0] shift_reg_out [0:SIZE-1]; // Shift register outputs

    // PWM module as clock divider for shift register
    pwm_module #(
        .bit_width(WIDTH)
    ) pwm_clk_div (
        .clk(clk),                      // Main clock
        .rst_n(rst_n),                  // Reset
        .duty(8'h80),                   // 50% duty cycle for slower clock
        .max_value(8'hFF),              // Full-range counter
        .pwm_out(slow_clk)              // PWM output used as shift register clock
    );

    // Shift register instance (uses PWM output as clock)
    shift_register #(
        .WIDTH(WIDTH),
        .SIZE(SIZE)
    ) shift_reg (
        .clk(gated_slow_clk),   // Slow PWM-generated clock
        .rst_n(rst_n),
        .data_in(ui_in),  // Inputs drive the shift register
        .reg_out(shift_reg_out)
    );

    // 8 PWM Modules, each fed by the shift register
    genvar i;
    generate
        for (i = 0; i < SIZE; i = i + 1) begin : pwm_gen
            pwm_module #(
                .bit_width(WIDTH)
            ) pwm_inst (
                .clk(clk),                      // PWM modules use main clock
                .rst_n(rst_n),                  // Reset
                .duty(shift_reg_out[i]),        // Shift register output as duty cycle
                .max_value(8'hFF),              // Max value = 255 (full range)
                .pwm_out(uo_out[i])             // PWM output mapped to `uo_out`
            );
        end
    endgenerate

    assign gated_slow_clk = (!rst_n) ? clk : slow_clk;

endmodule
